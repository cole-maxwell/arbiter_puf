* File: /home/ece658_2020/chmaxwell/lab5/part4/arbiter_puf.pex.netlist
* Created: Tue Dec  8 22:00:59 2020
* Program "Calibre xRC"
* Version "v2011.3_29.20"
* 


.include "/home/ece658_2020/chmaxwell/lab5/part4/arbiter_puf.pex.netlist.pex"
* include transistor models. include command can also be used to include other spice files
.include '$PDK_DIR/ncsu_basekit/models/hspice/hspice_nom.include'

* Analysis commands
.param vdd_val = 1.1
Vsupply vdd 0 vdd_val
Vgnd gnd 0 0

* Digital vector file for input from same directory
.vec 'arbiter_puf_input.vec'

* Simulation options
.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    POST

.subckt arbiter_puf  GND VDD Q_NOT Q R S SEL0 SEL1 SEL2 SEL3 SEL4 SEL5 SEL6 SEL7
* 
* SEL7	SEL7
* SEL6	SEL6
* SEL5	SEL5
* SEL4	SEL4
* SEL3	SEL3
* SEL2	SEL2
* SEL1	SEL1
* SEL0	SEL0
* S	S
* R	R
* Q	Q
* Q_NOT	Q_NOT
* VDD	VDD
* GND	GND
mXI8/MM0 N_Q_NOT_XI8/MM0_d N_NET32_XI8/MM0_g N_VDD_XI8/MM0_s N_VDD_XI8/MM0_b
+ PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI8/MM1 N_Q_NOT_XI8/MM0_d N_Q_XI8/MM1_g N_VDD_XI8/MM1_s N_VDD_XI8/MM0_b
+ PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI8/MM3 N_Q_XI8/MM3_d N_NET31_XI8/MM3_g N_VDD_XI8/MM3_s N_VDD_XI8/MM0_b
+ PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI8/MM2 N_Q_XI8/MM3_d N_Q_NOT_XI8/MM2_g N_VDD_XI8/MM2_s N_VDD_XI8/MM0_b
+ PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI8/MM5 XI8/NET24 N_NET32_XI8/MM5_g N_GND_XI8/MM5_s N_GND_XI8/MM5_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI8/MM4 N_Q_NOT_XI8/MM4_d N_Q_XI8/MM4_g XI8/NET24 N_GND_XI8/MM5_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI8/MM7 XI8/NET23 N_NET31_XI8/MM7_g N_GND_XI8/MM7_s N_GND_XI8/MM5_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI8/MM6 N_Q_XI8/MM6_d N_Q_NOT_XI8/MM6_g XI8/NET23 N_GND_XI8/MM5_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI6/XI6/MM0 N_XI6/NET19_XI6/XI6/MM0_d N_SEL0_XI6/XI6/MM0_g N_GND_XI6/XI6/MM0_s
+ N_GND_XI6/XI5/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI6/XI6/MM1 N_XI6/NET19_XI6/XI6/MM1_d N_SEL0_XI6/XI6/MM1_g N_VDD_XI6/XI6/MM1_s
+ N_VDD_XI6/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI6/XI1/MM2 N_XI6/NET22_XI6/XI1/MM2_d N_S_XI6/XI1/MM2_g N_VDD_XI6/XI1/MM2_s
+ N_VDD_XI6/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI1/MM3 N_XI6/NET22_XI6/XI1/MM2_d N_XI6/NET19_XI6/XI1/MM3_g
+ N_VDD_XI6/XI1/MM3_s N_VDD_XI6/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI6/XI5/MM2 N_XI6/NET25_XI6/XI5/MM2_d N_S_XI6/XI5/MM2_g N_VDD_XI6/XI5/MM2_s
+ N_VDD_XI6/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI5/MM3 N_XI6/NET25_XI6/XI5/MM2_d N_XI6/NET19_XI6/XI5/MM3_g
+ N_VDD_XI6/XI5/MM3_s N_VDD_XI6/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI6/XI0/MM2 N_XI6/NET24_XI6/XI0/MM2_d N_SEL0_XI6/XI0/MM2_g N_VDD_XI6/XI0/MM2_s
+ N_VDD_XI6/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI0/MM3 N_XI6/NET24_XI6/XI0/MM2_d N_R_XI6/XI0/MM3_g N_VDD_XI6/XI0/MM3_s
+ N_VDD_XI6/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI3/MM2 N_XI6/NET23_XI6/XI3/MM2_d N_SEL0_XI6/XI3/MM2_g N_VDD_XI6/XI3/MM2_s
+ N_VDD_XI6/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI3/MM3 N_XI6/NET23_XI6/XI3/MM2_d N_R_XI6/XI3/MM3_g N_VDD_XI6/XI3/MM3_s
+ N_VDD_XI6/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI2/MM2 N_NET46_XI6/XI2/MM2_d N_XI6/NET22_XI6/XI2/MM2_g N_VDD_XI6/XI2/MM2_s
+ N_VDD_XI6/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI2/MM3 N_NET46_XI6/XI2/MM2_d N_XI6/NET24_XI6/XI2/MM3_g N_VDD_XI6/XI2/MM3_s
+ N_VDD_XI6/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI4/MM3 N_NET45_XI6/XI4/MM3_d N_XI6/NET25_XI6/XI4/MM3_g N_VDD_XI6/XI4/MM3_s
+ N_VDD_XI6/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI4/MM2 N_NET45_XI6/XI4/MM3_d N_XI6/NET23_XI6/XI4/MM2_g N_VDD_XI6/XI4/MM2_s
+ N_VDD_XI6/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI1/MM1 XI6/XI1/NET16 N_S_XI6/XI1/MM1_g N_GND_XI6/XI1/MM1_s
+ N_GND_XI6/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI1/MM0 N_XI6/NET22_XI6/XI1/MM0_d N_XI6/NET19_XI6/XI1/MM0_g XI6/XI1/NET16
+ N_GND_XI6/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI6/XI5/MM1 XI6/XI5/NET16 N_S_XI6/XI5/MM1_g N_GND_XI6/XI5/MM1_s
+ N_GND_XI6/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI5/MM0 N_XI6/NET25_XI6/XI5/MM0_d N_XI6/NET19_XI6/XI5/MM0_g XI6/XI5/NET16
+ N_GND_XI6/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI6/XI0/MM1 XI6/XI0/NET16 N_SEL0_XI6/XI0/MM1_g N_GND_XI6/XI0/MM1_s
+ N_GND_XI6/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI0/MM0 N_XI6/NET24_XI6/XI0/MM0_d N_R_XI6/XI0/MM0_g XI6/XI0/NET16
+ N_GND_XI6/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI6/XI3/MM1 XI6/XI3/NET16 N_SEL0_XI6/XI3/MM1_g N_GND_XI6/XI3/MM1_s
+ N_GND_XI6/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI3/MM0 N_XI6/NET23_XI6/XI3/MM0_d N_R_XI6/XI3/MM0_g XI6/XI3/NET16
+ N_GND_XI6/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI6/XI2/MM1 XI6/XI2/NET16 N_XI6/NET22_XI6/XI2/MM1_g N_GND_XI6/XI2/MM1_s
+ N_GND_XI6/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI2/MM0 N_NET46_XI6/XI2/MM0_d N_XI6/NET24_XI6/XI2/MM0_g XI6/XI2/NET16
+ N_GND_XI6/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI6/XI4/MM0 XI6/XI4/NET16 N_XI6/NET25_XI6/XI4/MM0_g N_GND_XI6/XI4/MM0_s
+ N_GND_XI6/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI6/XI4/MM1 N_NET45_XI6/XI4/MM1_d N_XI6/NET23_XI6/XI4/MM1_g XI6/XI4/NET16
+ N_GND_XI6/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI6/MM0 N_XI2/NET19_XI2/XI6/MM0_d N_SEL1_XI2/XI6/MM0_g N_GND_XI2/XI6/MM0_s
+ N_GND_XI2/XI5/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI2/XI6/MM1 N_XI2/NET19_XI2/XI6/MM1_d N_SEL1_XI2/XI6/MM1_g N_VDD_XI2/XI6/MM1_s
+ N_VDD_XI2/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI2/XI1/MM2 N_XI2/NET22_XI2/XI1/MM2_d N_NET45_XI2/XI1/MM2_g N_VDD_XI2/XI1/MM2_s
+ N_VDD_XI2/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI1/MM3 N_XI2/NET22_XI2/XI1/MM2_d N_XI2/NET19_XI2/XI1/MM3_g
+ N_VDD_XI2/XI1/MM3_s N_VDD_XI2/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI2/XI5/MM2 N_XI2/NET25_XI2/XI5/MM2_d N_NET45_XI2/XI5/MM2_g N_VDD_XI2/XI5/MM2_s
+ N_VDD_XI2/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI5/MM3 N_XI2/NET25_XI2/XI5/MM2_d N_XI2/NET19_XI2/XI5/MM3_g
+ N_VDD_XI2/XI5/MM3_s N_VDD_XI2/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI2/XI0/MM2 N_XI2/NET24_XI2/XI0/MM2_d N_SEL1_XI2/XI0/MM2_g N_VDD_XI2/XI0/MM2_s
+ N_VDD_XI2/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI0/MM3 N_XI2/NET24_XI2/XI0/MM2_d N_NET46_XI2/XI0/MM3_g N_VDD_XI2/XI0/MM3_s
+ N_VDD_XI2/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI3/MM2 N_XI2/NET23_XI2/XI3/MM2_d N_SEL1_XI2/XI3/MM2_g N_VDD_XI2/XI3/MM2_s
+ N_VDD_XI2/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI3/MM3 N_XI2/NET23_XI2/XI3/MM2_d N_NET46_XI2/XI3/MM3_g N_VDD_XI2/XI3/MM3_s
+ N_VDD_XI2/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI2/MM2 N_NET44_XI2/XI2/MM2_d N_XI2/NET22_XI2/XI2/MM2_g N_VDD_XI2/XI2/MM2_s
+ N_VDD_XI2/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI2/MM3 N_NET44_XI2/XI2/MM2_d N_XI2/NET24_XI2/XI2/MM3_g N_VDD_XI2/XI2/MM3_s
+ N_VDD_XI2/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI4/MM3 N_NET43_XI2/XI4/MM3_d N_XI2/NET25_XI2/XI4/MM3_g N_VDD_XI2/XI4/MM3_s
+ N_VDD_XI2/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI4/MM2 N_NET43_XI2/XI4/MM3_d N_XI2/NET23_XI2/XI4/MM2_g N_VDD_XI2/XI4/MM2_s
+ N_VDD_XI2/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI1/MM1 XI2/XI1/NET16 N_NET45_XI2/XI1/MM1_g N_GND_XI2/XI1/MM1_s
+ N_GND_XI2/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI1/MM0 N_XI2/NET22_XI2/XI1/MM0_d N_XI2/NET19_XI2/XI1/MM0_g XI2/XI1/NET16
+ N_GND_XI2/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI5/MM1 XI2/XI5/NET16 N_NET45_XI2/XI5/MM1_g N_GND_XI2/XI5/MM1_s
+ N_GND_XI2/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI5/MM0 N_XI2/NET25_XI2/XI5/MM0_d N_XI2/NET19_XI2/XI5/MM0_g XI2/XI5/NET16
+ N_GND_XI2/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI0/MM1 XI2/XI0/NET16 N_SEL1_XI2/XI0/MM1_g N_GND_XI2/XI0/MM1_s
+ N_GND_XI2/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI0/MM0 N_XI2/NET24_XI2/XI0/MM0_d N_NET46_XI2/XI0/MM0_g XI2/XI0/NET16
+ N_GND_XI2/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI3/MM1 XI2/XI3/NET16 N_SEL1_XI2/XI3/MM1_g N_GND_XI2/XI3/MM1_s
+ N_GND_XI2/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI3/MM0 N_XI2/NET23_XI2/XI3/MM0_d N_NET46_XI2/XI3/MM0_g XI2/XI3/NET16
+ N_GND_XI2/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI2/MM1 XI2/XI2/NET16 N_XI2/NET22_XI2/XI2/MM1_g N_GND_XI2/XI2/MM1_s
+ N_GND_XI2/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI2/MM0 N_NET44_XI2/XI2/MM0_d N_XI2/NET24_XI2/XI2/MM0_g XI2/XI2/NET16
+ N_GND_XI2/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI4/MM0 XI2/XI4/NET16 N_XI2/NET25_XI2/XI4/MM0_g N_GND_XI2/XI4/MM0_s
+ N_GND_XI2/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI4/MM1 N_NET43_XI2/XI4/MM1_d N_XI2/NET23_XI2/XI4/MM1_g XI2/XI4/NET16
+ N_GND_XI2/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI6/MM0 N_XI1/NET19_XI1/XI6/MM0_d N_SEL2_XI1/XI6/MM0_g N_GND_XI1/XI6/MM0_s
+ N_GND_XI1/XI5/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI1/XI6/MM1 N_XI1/NET19_XI1/XI6/MM1_d N_SEL2_XI1/XI6/MM1_g N_VDD_XI1/XI6/MM1_s
+ N_VDD_XI1/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI1/XI1/MM2 N_XI1/NET22_XI1/XI1/MM2_d N_NET43_XI1/XI1/MM2_g N_VDD_XI1/XI1/MM2_s
+ N_VDD_XI1/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI1/MM3 N_XI1/NET22_XI1/XI1/MM2_d N_XI1/NET19_XI1/XI1/MM3_g
+ N_VDD_XI1/XI1/MM3_s N_VDD_XI1/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI1/XI5/MM2 N_XI1/NET25_XI1/XI5/MM2_d N_NET43_XI1/XI5/MM2_g N_VDD_XI1/XI5/MM2_s
+ N_VDD_XI1/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI5/MM3 N_XI1/NET25_XI1/XI5/MM2_d N_XI1/NET19_XI1/XI5/MM3_g
+ N_VDD_XI1/XI5/MM3_s N_VDD_XI1/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI1/XI0/MM2 N_XI1/NET24_XI1/XI0/MM2_d N_SEL2_XI1/XI0/MM2_g N_VDD_XI1/XI0/MM2_s
+ N_VDD_XI1/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI0/MM3 N_XI1/NET24_XI1/XI0/MM2_d N_NET44_XI1/XI0/MM3_g N_VDD_XI1/XI0/MM3_s
+ N_VDD_XI1/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI3/MM2 N_XI1/NET23_XI1/XI3/MM2_d N_SEL2_XI1/XI3/MM2_g N_VDD_XI1/XI3/MM2_s
+ N_VDD_XI1/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI3/MM3 N_XI1/NET23_XI1/XI3/MM2_d N_NET44_XI1/XI3/MM3_g N_VDD_XI1/XI3/MM3_s
+ N_VDD_XI1/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI2/MM2 N_NET42_XI1/XI2/MM2_d N_XI1/NET22_XI1/XI2/MM2_g N_VDD_XI1/XI2/MM2_s
+ N_VDD_XI1/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI2/MM3 N_NET42_XI1/XI2/MM2_d N_XI1/NET24_XI1/XI2/MM3_g N_VDD_XI1/XI2/MM3_s
+ N_VDD_XI1/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI4/MM3 N_NET41_XI1/XI4/MM3_d N_XI1/NET25_XI1/XI4/MM3_g N_VDD_XI1/XI4/MM3_s
+ N_VDD_XI1/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI4/MM2 N_NET41_XI1/XI4/MM3_d N_XI1/NET23_XI1/XI4/MM2_g N_VDD_XI1/XI4/MM2_s
+ N_VDD_XI1/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI1/MM1 XI1/XI1/NET16 N_NET43_XI1/XI1/MM1_g N_GND_XI1/XI1/MM1_s
+ N_GND_XI1/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI1/MM0 N_XI1/NET22_XI1/XI1/MM0_d N_XI1/NET19_XI1/XI1/MM0_g XI1/XI1/NET16
+ N_GND_XI1/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI5/MM1 XI1/XI5/NET16 N_NET43_XI1/XI5/MM1_g N_GND_XI1/XI5/MM1_s
+ N_GND_XI1/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI5/MM0 N_XI1/NET25_XI1/XI5/MM0_d N_XI1/NET19_XI1/XI5/MM0_g XI1/XI5/NET16
+ N_GND_XI1/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI0/MM1 XI1/XI0/NET16 N_SEL2_XI1/XI0/MM1_g N_GND_XI1/XI0/MM1_s
+ N_GND_XI1/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI0/MM0 N_XI1/NET24_XI1/XI0/MM0_d N_NET44_XI1/XI0/MM0_g XI1/XI0/NET16
+ N_GND_XI1/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI3/MM1 XI1/XI3/NET16 N_SEL2_XI1/XI3/MM1_g N_GND_XI1/XI3/MM1_s
+ N_GND_XI1/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI3/MM0 N_XI1/NET23_XI1/XI3/MM0_d N_NET44_XI1/XI3/MM0_g XI1/XI3/NET16
+ N_GND_XI1/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI2/MM1 XI1/XI2/NET16 N_XI1/NET22_XI1/XI2/MM1_g N_GND_XI1/XI2/MM1_s
+ N_GND_XI1/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI2/MM0 N_NET42_XI1/XI2/MM0_d N_XI1/NET24_XI1/XI2/MM0_g XI1/XI2/NET16
+ N_GND_XI1/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI4/MM0 XI1/XI4/NET16 N_XI1/NET25_XI1/XI4/MM0_g N_GND_XI1/XI4/MM0_s
+ N_GND_XI1/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI4/MM1 N_NET41_XI1/XI4/MM1_d N_XI1/NET23_XI1/XI4/MM1_g XI1/XI4/NET16
+ N_GND_XI1/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI0/XI6/MM0 N_XI0/NET19_XI0/XI6/MM0_d N_SEL3_XI0/XI6/MM0_g N_GND_XI0/XI6/MM0_s
+ N_GND_XI0/XI5/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI0/XI6/MM1 N_XI0/NET19_XI0/XI6/MM1_d N_SEL3_XI0/XI6/MM1_g N_VDD_XI0/XI6/MM1_s
+ N_VDD_XI0/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI0/XI1/MM2 N_XI0/NET22_XI0/XI1/MM2_d N_NET41_XI0/XI1/MM2_g N_VDD_XI0/XI1/MM2_s
+ N_VDD_XI0/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI1/MM3 N_XI0/NET22_XI0/XI1/MM2_d N_XI0/NET19_XI0/XI1/MM3_g
+ N_VDD_XI0/XI1/MM3_s N_VDD_XI0/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI0/XI5/MM2 N_XI0/NET25_XI0/XI5/MM2_d N_NET41_XI0/XI5/MM2_g N_VDD_XI0/XI5/MM2_s
+ N_VDD_XI0/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI5/MM3 N_XI0/NET25_XI0/XI5/MM2_d N_XI0/NET19_XI0/XI5/MM3_g
+ N_VDD_XI0/XI5/MM3_s N_VDD_XI0/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI0/XI0/MM2 N_XI0/NET24_XI0/XI0/MM2_d N_SEL3_XI0/XI0/MM2_g N_VDD_XI0/XI0/MM2_s
+ N_VDD_XI0/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI0/MM3 N_XI0/NET24_XI0/XI0/MM2_d N_NET42_XI0/XI0/MM3_g N_VDD_XI0/XI0/MM3_s
+ N_VDD_XI0/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI3/MM2 N_XI0/NET23_XI0/XI3/MM2_d N_SEL3_XI0/XI3/MM2_g N_VDD_XI0/XI3/MM2_s
+ N_VDD_XI0/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI3/MM3 N_XI0/NET23_XI0/XI3/MM2_d N_NET42_XI0/XI3/MM3_g N_VDD_XI0/XI3/MM3_s
+ N_VDD_XI0/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI2/MM2 N_NET40_XI0/XI2/MM2_d N_XI0/NET22_XI0/XI2/MM2_g N_VDD_XI0/XI2/MM2_s
+ N_VDD_XI0/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI2/MM3 N_NET40_XI0/XI2/MM2_d N_XI0/NET24_XI0/XI2/MM3_g N_VDD_XI0/XI2/MM3_s
+ N_VDD_XI0/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI4/MM3 N_NET39_XI0/XI4/MM3_d N_XI0/NET25_XI0/XI4/MM3_g N_VDD_XI0/XI4/MM3_s
+ N_VDD_XI0/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI4/MM2 N_NET39_XI0/XI4/MM3_d N_XI0/NET23_XI0/XI4/MM2_g N_VDD_XI0/XI4/MM2_s
+ N_VDD_XI0/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI1/MM1 XI0/XI1/NET16 N_NET41_XI0/XI1/MM1_g N_GND_XI0/XI1/MM1_s
+ N_GND_XI0/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI1/MM0 N_XI0/NET22_XI0/XI1/MM0_d N_XI0/NET19_XI0/XI1/MM0_g XI0/XI1/NET16
+ N_GND_XI0/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI0/XI5/MM1 XI0/XI5/NET16 N_NET41_XI0/XI5/MM1_g N_GND_XI0/XI5/MM1_s
+ N_GND_XI0/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI5/MM0 N_XI0/NET25_XI0/XI5/MM0_d N_XI0/NET19_XI0/XI5/MM0_g XI0/XI5/NET16
+ N_GND_XI0/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI0/XI0/MM1 XI0/XI0/NET16 N_SEL3_XI0/XI0/MM1_g N_GND_XI0/XI0/MM1_s
+ N_GND_XI0/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI0/MM0 N_XI0/NET24_XI0/XI0/MM0_d N_NET42_XI0/XI0/MM0_g XI0/XI0/NET16
+ N_GND_XI0/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI0/XI3/MM1 XI0/XI3/NET16 N_SEL3_XI0/XI3/MM1_g N_GND_XI0/XI3/MM1_s
+ N_GND_XI0/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI3/MM0 N_XI0/NET23_XI0/XI3/MM0_d N_NET42_XI0/XI3/MM0_g XI0/XI3/NET16
+ N_GND_XI0/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI0/XI2/MM1 XI0/XI2/NET16 N_XI0/NET22_XI0/XI2/MM1_g N_GND_XI0/XI2/MM1_s
+ N_GND_XI0/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI2/MM0 N_NET40_XI0/XI2/MM0_d N_XI0/NET24_XI0/XI2/MM0_g XI0/XI2/NET16
+ N_GND_XI0/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI0/XI4/MM0 XI0/XI4/NET16 N_XI0/NET25_XI0/XI4/MM0_g N_GND_XI0/XI4/MM0_s
+ N_GND_XI0/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI4/MM1 N_NET39_XI0/XI4/MM1_d N_XI0/NET23_XI0/XI4/MM1_g XI0/XI4/NET16
+ N_GND_XI0/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI6/MM0 N_XI3/NET19_XI3/XI6/MM0_d N_SEL4_XI3/XI6/MM0_g N_GND_XI3/XI6/MM0_s
+ N_GND_XI3/XI5/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI3/XI6/MM1 N_XI3/NET19_XI3/XI6/MM1_d N_SEL4_XI3/XI6/MM1_g N_VDD_XI3/XI6/MM1_s
+ N_VDD_XI3/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI3/XI1/MM2 N_XI3/NET22_XI3/XI1/MM2_d N_NET39_XI3/XI1/MM2_g N_VDD_XI3/XI1/MM2_s
+ N_VDD_XI3/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI1/MM3 N_XI3/NET22_XI3/XI1/MM2_d N_XI3/NET19_XI3/XI1/MM3_g
+ N_VDD_XI3/XI1/MM3_s N_VDD_XI3/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI3/XI5/MM2 N_XI3/NET25_XI3/XI5/MM2_d N_NET39_XI3/XI5/MM2_g N_VDD_XI3/XI5/MM2_s
+ N_VDD_XI3/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI5/MM3 N_XI3/NET25_XI3/XI5/MM2_d N_XI3/NET19_XI3/XI5/MM3_g
+ N_VDD_XI3/XI5/MM3_s N_VDD_XI3/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI3/XI0/MM2 N_XI3/NET24_XI3/XI0/MM2_d N_SEL4_XI3/XI0/MM2_g N_VDD_XI3/XI0/MM2_s
+ N_VDD_XI3/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI0/MM3 N_XI3/NET24_XI3/XI0/MM2_d N_NET40_XI3/XI0/MM3_g N_VDD_XI3/XI0/MM3_s
+ N_VDD_XI3/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI3/MM2 N_XI3/NET23_XI3/XI3/MM2_d N_SEL4_XI3/XI3/MM2_g N_VDD_XI3/XI3/MM2_s
+ N_VDD_XI3/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI3/MM3 N_XI3/NET23_XI3/XI3/MM2_d N_NET40_XI3/XI3/MM3_g N_VDD_XI3/XI3/MM3_s
+ N_VDD_XI3/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI2/MM2 N_NET38_XI3/XI2/MM2_d N_XI3/NET22_XI3/XI2/MM2_g N_VDD_XI3/XI2/MM2_s
+ N_VDD_XI3/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI2/MM3 N_NET38_XI3/XI2/MM2_d N_XI3/NET24_XI3/XI2/MM3_g N_VDD_XI3/XI2/MM3_s
+ N_VDD_XI3/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI4/MM3 N_NET37_XI3/XI4/MM3_d N_XI3/NET25_XI3/XI4/MM3_g N_VDD_XI3/XI4/MM3_s
+ N_VDD_XI3/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI4/MM2 N_NET37_XI3/XI4/MM3_d N_XI3/NET23_XI3/XI4/MM2_g N_VDD_XI3/XI4/MM2_s
+ N_VDD_XI3/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI1/MM1 XI3/XI1/NET16 N_NET39_XI3/XI1/MM1_g N_GND_XI3/XI1/MM1_s
+ N_GND_XI3/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI1/MM0 N_XI3/NET22_XI3/XI1/MM0_d N_XI3/NET19_XI3/XI1/MM0_g XI3/XI1/NET16
+ N_GND_XI3/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI5/MM1 XI3/XI5/NET16 N_NET39_XI3/XI5/MM1_g N_GND_XI3/XI5/MM1_s
+ N_GND_XI3/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI5/MM0 N_XI3/NET25_XI3/XI5/MM0_d N_XI3/NET19_XI3/XI5/MM0_g XI3/XI5/NET16
+ N_GND_XI3/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI0/MM1 XI3/XI0/NET16 N_SEL4_XI3/XI0/MM1_g N_GND_XI3/XI0/MM1_s
+ N_GND_XI3/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI0/MM0 N_XI3/NET24_XI3/XI0/MM0_d N_NET40_XI3/XI0/MM0_g XI3/XI0/NET16
+ N_GND_XI3/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI3/MM1 XI3/XI3/NET16 N_SEL4_XI3/XI3/MM1_g N_GND_XI3/XI3/MM1_s
+ N_GND_XI3/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI3/MM0 N_XI3/NET23_XI3/XI3/MM0_d N_NET40_XI3/XI3/MM0_g XI3/XI3/NET16
+ N_GND_XI3/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI2/MM1 XI3/XI2/NET16 N_XI3/NET22_XI3/XI2/MM1_g N_GND_XI3/XI2/MM1_s
+ N_GND_XI3/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI2/MM0 N_NET38_XI3/XI2/MM0_d N_XI3/NET24_XI3/XI2/MM0_g XI3/XI2/NET16
+ N_GND_XI3/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI4/MM0 XI3/XI4/NET16 N_XI3/NET25_XI3/XI4/MM0_g N_GND_XI3/XI4/MM0_s
+ N_GND_XI3/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI4/MM1 N_NET37_XI3/XI4/MM1_d N_XI3/NET23_XI3/XI4/MM1_g XI3/XI4/NET16
+ N_GND_XI3/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI4/XI6/MM0 N_XI4/NET19_XI4/XI6/MM0_d N_SEL5_XI4/XI6/MM0_g N_GND_XI4/XI6/MM0_s
+ N_GND_XI4/XI5/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI4/XI6/MM1 N_XI4/NET19_XI4/XI6/MM1_d N_SEL5_XI4/XI6/MM1_g N_VDD_XI4/XI6/MM1_s
+ N_VDD_XI4/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI4/XI1/MM2 N_XI4/NET22_XI4/XI1/MM2_d N_NET37_XI4/XI1/MM2_g N_VDD_XI4/XI1/MM2_s
+ N_VDD_XI4/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI1/MM3 N_XI4/NET22_XI4/XI1/MM2_d N_XI4/NET19_XI4/XI1/MM3_g
+ N_VDD_XI4/XI1/MM3_s N_VDD_XI4/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI4/XI5/MM2 N_XI4/NET25_XI4/XI5/MM2_d N_NET37_XI4/XI5/MM2_g N_VDD_XI4/XI5/MM2_s
+ N_VDD_XI4/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI5/MM3 N_XI4/NET25_XI4/XI5/MM2_d N_XI4/NET19_XI4/XI5/MM3_g
+ N_VDD_XI4/XI5/MM3_s N_VDD_XI4/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI4/XI0/MM2 N_XI4/NET24_XI4/XI0/MM2_d N_SEL5_XI4/XI0/MM2_g N_VDD_XI4/XI0/MM2_s
+ N_VDD_XI4/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI0/MM3 N_XI4/NET24_XI4/XI0/MM2_d N_NET38_XI4/XI0/MM3_g N_VDD_XI4/XI0/MM3_s
+ N_VDD_XI4/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI3/MM2 N_XI4/NET23_XI4/XI3/MM2_d N_SEL5_XI4/XI3/MM2_g N_VDD_XI4/XI3/MM2_s
+ N_VDD_XI4/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI3/MM3 N_XI4/NET23_XI4/XI3/MM2_d N_NET38_XI4/XI3/MM3_g N_VDD_XI4/XI3/MM3_s
+ N_VDD_XI4/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI2/MM2 N_NET36_XI4/XI2/MM2_d N_XI4/NET22_XI4/XI2/MM2_g N_VDD_XI4/XI2/MM2_s
+ N_VDD_XI4/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI2/MM3 N_NET36_XI4/XI2/MM2_d N_XI4/NET24_XI4/XI2/MM3_g N_VDD_XI4/XI2/MM3_s
+ N_VDD_XI4/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI4/MM3 N_NET35_XI4/XI4/MM3_d N_XI4/NET25_XI4/XI4/MM3_g N_VDD_XI4/XI4/MM3_s
+ N_VDD_XI4/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI4/MM2 N_NET35_XI4/XI4/MM3_d N_XI4/NET23_XI4/XI4/MM2_g N_VDD_XI4/XI4/MM2_s
+ N_VDD_XI4/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI1/MM1 XI4/XI1/NET16 N_NET37_XI4/XI1/MM1_g N_GND_XI4/XI1/MM1_s
+ N_GND_XI4/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI1/MM0 N_XI4/NET22_XI4/XI1/MM0_d N_XI4/NET19_XI4/XI1/MM0_g XI4/XI1/NET16
+ N_GND_XI4/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI4/XI5/MM1 XI4/XI5/NET16 N_NET37_XI4/XI5/MM1_g N_GND_XI4/XI5/MM1_s
+ N_GND_XI4/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI5/MM0 N_XI4/NET25_XI4/XI5/MM0_d N_XI4/NET19_XI4/XI5/MM0_g XI4/XI5/NET16
+ N_GND_XI4/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI4/XI0/MM1 XI4/XI0/NET16 N_SEL5_XI4/XI0/MM1_g N_GND_XI4/XI0/MM1_s
+ N_GND_XI4/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI0/MM0 N_XI4/NET24_XI4/XI0/MM0_d N_NET38_XI4/XI0/MM0_g XI4/XI0/NET16
+ N_GND_XI4/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI4/XI3/MM1 XI4/XI3/NET16 N_SEL5_XI4/XI3/MM1_g N_GND_XI4/XI3/MM1_s
+ N_GND_XI4/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI3/MM0 N_XI4/NET23_XI4/XI3/MM0_d N_NET38_XI4/XI3/MM0_g XI4/XI3/NET16
+ N_GND_XI4/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI4/XI2/MM1 XI4/XI2/NET16 N_XI4/NET22_XI4/XI2/MM1_g N_GND_XI4/XI2/MM1_s
+ N_GND_XI4/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI2/MM0 N_NET36_XI4/XI2/MM0_d N_XI4/NET24_XI4/XI2/MM0_g XI4/XI2/NET16
+ N_GND_XI4/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI4/XI4/MM0 XI4/XI4/NET16 N_XI4/NET25_XI4/XI4/MM0_g N_GND_XI4/XI4/MM0_s
+ N_GND_XI4/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI4/XI4/MM1 N_NET35_XI4/XI4/MM1_d N_XI4/NET23_XI4/XI4/MM1_g XI4/XI4/NET16
+ N_GND_XI4/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI5/XI6/MM0 N_XI5/NET19_XI5/XI6/MM0_d N_SEL6_XI5/XI6/MM0_g N_GND_XI5/XI6/MM0_s
+ N_GND_XI5/XI5/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI5/XI6/MM1 N_XI5/NET19_XI5/XI6/MM1_d N_SEL6_XI5/XI6/MM1_g N_VDD_XI5/XI6/MM1_s
+ N_VDD_XI5/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI5/XI1/MM2 N_XI5/NET22_XI5/XI1/MM2_d N_NET35_XI5/XI1/MM2_g N_VDD_XI5/XI1/MM2_s
+ N_VDD_XI5/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI1/MM3 N_XI5/NET22_XI5/XI1/MM2_d N_XI5/NET19_XI5/XI1/MM3_g
+ N_VDD_XI5/XI1/MM3_s N_VDD_XI5/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI5/XI5/MM2 N_XI5/NET25_XI5/XI5/MM2_d N_NET35_XI5/XI5/MM2_g N_VDD_XI5/XI5/MM2_s
+ N_VDD_XI5/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI5/MM3 N_XI5/NET25_XI5/XI5/MM2_d N_XI5/NET19_XI5/XI5/MM3_g
+ N_VDD_XI5/XI5/MM3_s N_VDD_XI5/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI5/XI0/MM2 N_XI5/NET24_XI5/XI0/MM2_d N_SEL6_XI5/XI0/MM2_g N_VDD_XI5/XI0/MM2_s
+ N_VDD_XI5/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI0/MM3 N_XI5/NET24_XI5/XI0/MM2_d N_NET36_XI5/XI0/MM3_g N_VDD_XI5/XI0/MM3_s
+ N_VDD_XI5/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI3/MM2 N_XI5/NET23_XI5/XI3/MM2_d N_SEL6_XI5/XI3/MM2_g N_VDD_XI5/XI3/MM2_s
+ N_VDD_XI5/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI3/MM3 N_XI5/NET23_XI5/XI3/MM2_d N_NET36_XI5/XI3/MM3_g N_VDD_XI5/XI3/MM3_s
+ N_VDD_XI5/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI2/MM2 N_NET34_XI5/XI2/MM2_d N_XI5/NET22_XI5/XI2/MM2_g N_VDD_XI5/XI2/MM2_s
+ N_VDD_XI5/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI2/MM3 N_NET34_XI5/XI2/MM2_d N_XI5/NET24_XI5/XI2/MM3_g N_VDD_XI5/XI2/MM3_s
+ N_VDD_XI5/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI4/MM3 N_NET33_XI5/XI4/MM3_d N_XI5/NET25_XI5/XI4/MM3_g N_VDD_XI5/XI4/MM3_s
+ N_VDD_XI5/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI4/MM2 N_NET33_XI5/XI4/MM3_d N_XI5/NET23_XI5/XI4/MM2_g N_VDD_XI5/XI4/MM2_s
+ N_VDD_XI5/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI1/MM1 XI5/XI1/NET16 N_NET35_XI5/XI1/MM1_g N_GND_XI5/XI1/MM1_s
+ N_GND_XI5/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI1/MM0 N_XI5/NET22_XI5/XI1/MM0_d N_XI5/NET19_XI5/XI1/MM0_g XI5/XI1/NET16
+ N_GND_XI5/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI5/XI5/MM1 XI5/XI5/NET16 N_NET35_XI5/XI5/MM1_g N_GND_XI5/XI5/MM1_s
+ N_GND_XI5/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI5/MM0 N_XI5/NET25_XI5/XI5/MM0_d N_XI5/NET19_XI5/XI5/MM0_g XI5/XI5/NET16
+ N_GND_XI5/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI5/XI0/MM1 XI5/XI0/NET16 N_SEL6_XI5/XI0/MM1_g N_GND_XI5/XI0/MM1_s
+ N_GND_XI5/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI0/MM0 N_XI5/NET24_XI5/XI0/MM0_d N_NET36_XI5/XI0/MM0_g XI5/XI0/NET16
+ N_GND_XI5/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI5/XI3/MM1 XI5/XI3/NET16 N_SEL6_XI5/XI3/MM1_g N_GND_XI5/XI3/MM1_s
+ N_GND_XI5/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI3/MM0 N_XI5/NET23_XI5/XI3/MM0_d N_NET36_XI5/XI3/MM0_g XI5/XI3/NET16
+ N_GND_XI5/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI5/XI2/MM1 XI5/XI2/NET16 N_XI5/NET22_XI5/XI2/MM1_g N_GND_XI5/XI2/MM1_s
+ N_GND_XI5/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI2/MM0 N_NET34_XI5/XI2/MM0_d N_XI5/NET24_XI5/XI2/MM0_g XI5/XI2/NET16
+ N_GND_XI5/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI5/XI4/MM0 XI5/XI4/NET16 N_XI5/NET25_XI5/XI4/MM0_g N_GND_XI5/XI4/MM0_s
+ N_GND_XI5/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI5/XI4/MM1 N_NET33_XI5/XI4/MM1_d N_XI5/NET23_XI5/XI4/MM1_g XI5/XI4/NET16
+ N_GND_XI5/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI7/XI6/MM0 N_XI7/NET19_XI7/XI6/MM0_d N_SEL7_XI7/XI6/MM0_g N_GND_XI7/XI6/MM0_s
+ N_GND_XI7/XI1/MM1_b NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15
+ PD=3.9e-07 PS=3.9e-07
mXI7/XI6/MM1 N_XI7/NET19_XI7/XI6/MM1_d N_SEL7_XI7/XI6/MM1_g N_VDD_XI7/XI6/MM1_s
+ N_VDD_XI7/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14
+ PD=5.7e-07 PS=5.7e-07
mXI7/XI5/MM2 N_XI7/NET25_XI7/XI5/MM2_d N_NET33_XI7/XI5/MM2_g N_VDD_XI7/XI5/MM2_s
+ N_VDD_XI7/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI5/MM3 N_XI7/NET25_XI7/XI5/MM2_d N_XI7/NET19_XI7/XI5/MM3_g
+ N_VDD_XI7/XI5/MM3_s N_VDD_XI7/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI7/XI1/MM2 N_XI7/NET22_XI7/XI1/MM2_d N_NET33_XI7/XI1/MM2_g N_VDD_XI7/XI1/MM2_s
+ N_VDD_XI7/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI1/MM3 N_XI7/NET22_XI7/XI1/MM2_d N_XI7/NET19_XI7/XI1/MM3_g
+ N_VDD_XI7/XI1/MM3_s N_VDD_XI7/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14
+ AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI7/XI3/MM2 N_XI7/NET23_XI7/XI3/MM2_d N_SEL7_XI7/XI3/MM2_g N_VDD_XI7/XI3/MM2_s
+ N_VDD_XI7/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI3/MM3 N_XI7/NET23_XI7/XI3/MM2_d N_NET34_XI7/XI3/MM3_g N_VDD_XI7/XI3/MM3_s
+ N_VDD_XI7/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI0/MM2 N_XI7/NET24_XI7/XI0/MM2_d N_SEL7_XI7/XI0/MM2_g N_VDD_XI7/XI0/MM2_s
+ N_VDD_XI7/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI0/MM3 N_XI7/NET24_XI7/XI0/MM2_d N_NET34_XI7/XI0/MM3_g N_VDD_XI7/XI0/MM3_s
+ N_VDD_XI7/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI4/MM3 N_NET31_XI7/XI4/MM3_d N_XI7/NET25_XI7/XI4/MM3_g N_VDD_XI7/XI4/MM3_s
+ N_VDD_XI7/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI4/MM2 N_NET31_XI7/XI4/MM3_d N_XI7/NET23_XI7/XI4/MM2_g N_VDD_XI7/XI4/MM2_s
+ N_VDD_XI7/XI5/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI2/MM2 N_NET32_XI7/XI2/MM2_d N_XI7/NET22_XI7/XI2/MM2_g N_VDD_XI7/XI2/MM2_s
+ N_VDD_XI7/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI2/MM3 N_NET32_XI7/XI2/MM2_d N_XI7/NET24_XI7/XI2/MM3_g N_VDD_XI7/XI2/MM3_s
+ N_VDD_XI7/XI1/MM2_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI5/MM1 XI7/XI5/NET16 N_NET33_XI7/XI5/MM1_g N_GND_XI7/XI5/MM1_s
+ N_GND_XI7/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI5/MM0 N_XI7/NET25_XI7/XI5/MM0_d N_XI7/NET19_XI7/XI5/MM0_g XI7/XI5/NET16
+ N_GND_XI7/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI7/XI1/MM1 XI7/XI1/NET16 N_NET33_XI7/XI1/MM1_g N_GND_XI7/XI1/MM1_s
+ N_GND_XI7/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI1/MM0 N_XI7/NET22_XI7/XI1/MM0_d N_XI7/NET19_XI7/XI1/MM0_g XI7/XI1/NET16
+ N_GND_XI7/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI7/XI3/MM1 XI7/XI3/NET16 N_SEL7_XI7/XI3/MM1_g N_GND_XI7/XI3/MM1_s
+ N_GND_XI7/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI3/MM0 N_XI7/NET23_XI7/XI3/MM0_d N_NET34_XI7/XI3/MM0_g XI7/XI3/NET16
+ N_GND_XI7/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI7/XI0/MM1 XI7/XI0/NET16 N_SEL7_XI7/XI0/MM1_g N_GND_XI7/XI0/MM1_s
+ N_GND_XI7/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI0/MM0 N_XI7/NET24_XI7/XI0/MM0_d N_NET34_XI7/XI0/MM0_g XI7/XI0/NET16
+ N_GND_XI7/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI7/XI4/MM0 XI7/XI4/NET16 N_XI7/NET25_XI7/XI4/MM0_g N_GND_XI7/XI4/MM0_s
+ N_GND_XI7/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI4/MM1 N_NET31_XI7/XI4/MM1_d N_XI7/NET23_XI7/XI4/MM1_g XI7/XI4/NET16
+ N_GND_XI7/XI5/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI7/XI2/MM1 XI7/XI2/NET16 N_XI7/NET22_XI7/XI2/MM1_g N_GND_XI7/XI2/MM1_s
+ N_GND_XI7/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI7/XI2/MM0 N_NET32_XI7/XI2/MM0_d N_XI7/NET24_XI7/XI2/MM0_g XI7/XI2/NET16
+ N_GND_XI7/XI1/MM1_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
*
.include "/home/ece658_2020/chmaxwell/lab5/part4/arbiter_puf.pex.netlist.ARBITER_PUF.pxi"
*
.ends
*
*
x1 GND VDD Q_NOT Q R S SEL0 SEL1 SEL2 SEL3 SEL4 SEL5 SEL6 SEL7 ARBITER_PUF

*------------------------------------------------------------------------
* Stimulus
*------------------------------------------------------------------------

.tran 1p 600p

.END
